module sumador (
	input clk, rst,
   input [9:0] switches,
	output suma
);

suma_anterior	

endmodule